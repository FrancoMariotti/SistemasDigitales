library IEEE;
use IEEE.std_logic_1164.all;

entity mux4b is

end;


architecture mux4b_arq of mux4b is
	--parte declarativa
begin
	--parte descriptiva
end mux4b_arq;
